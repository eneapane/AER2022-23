package AcceleratorChecker;
    import MyTypes::*;
    import GetPut::*;
    import ClientServer::*;
    import FIFO::*;
    import ImageFunctions::*;
    import Gauss::*;
    import StmtFSM::*;
    import Settings::*;
    import Vector::*;
    import Top::*;

    module mkAcceleratorChecker(Empty);
        // TODO: Task 4.4
    endmodule
endpackage : AcceleratorChecker