package BufferTb;
    import MyTypes::*;
    import Settings::*;
    import Buffer::*;
    import FIFO::*;
    import GetPut::*;
    import ClientServer::*;
    import StmtFSM::*;

    module mkBufferTb(Empty);
        // TODO: Implement this module (task 3.1e)

    endmodule : mkBufferTb


endpackage : BufferTb