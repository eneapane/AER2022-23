package Settings;
  Integer width = 1173;
  Integer height = 470;
  Integer n_vals = width * height;
endpackage