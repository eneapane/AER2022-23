package Settings;
  // TODO: change width and height to fit your input image
  Integer width = 1173;
  Integer height = 470;
  Integer n_vals = width * height;

endpackage