package MyTypes;

typedef Bit#(8) GrayScale;

endpackage
