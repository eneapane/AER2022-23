package GaussChecker;
    import MyTypes::*;
    import GetPut::*;
    import ClientServer::*;
    import FIFO::*;
    import ImageFunctions::*;
    import Gauss::*;
    import StmtFSM::*;
    import Settings::*;
    import Vector::*;

    module mkGaussChecker(Empty);
        // TODO: implement me (task 3.1c)
    endmodule : mkGaussChecker
endpackage : GaussChecker